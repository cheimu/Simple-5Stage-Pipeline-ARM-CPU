module RegisterFile();

endmodule
